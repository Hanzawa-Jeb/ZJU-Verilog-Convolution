`ifdef VERILATE
    localparam DATA_FILE_PATH = "initial_data.hex";
`else
    localparam DATA_FILE_PATH = // fill the path;
`endif