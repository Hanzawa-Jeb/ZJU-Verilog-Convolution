`ifdef VERILATE
    localparam DATA_FILE_PATH = "initial_data.hex";
`else
    localparam DATA_FILE_PATH = "D:\\sysI\\sys1-sp25\\repo\\sys-project\\lab4-1\\syn\\initial_data.hex";
`endif